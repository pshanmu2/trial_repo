module my_verilog();

  //Preethi - TODO - Add my verilog code here later
endmodule
